

SAUS2US3US4US5US6US7US8US9US0USJU
DAUD2UD3UD4UD5UD6UD7UD8UD9UD0U
CAUC2UC3UC4UC5UC6UC7UC8UC9UC0U
HAUH2UH3UH4UH5UH6UH7UH8UH9UH0UHJU

CKUHQU
HKUCQU
SKUDQUCJU
DKUSQUDJU


